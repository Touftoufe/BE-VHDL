-- SoC.vhd

-- Generated using ACDS version 18.1 625

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity SoC is
	port (
		anemometer_data_anemometre_new_signal    : out std_logic_vector(7 downto 0);                    --    anemometer_data_anemometre.new_signal
		anemometer_data_valid_new_signal         : out std_logic;                                       --         anemometer_data_valid.new_signal
		anemometer_in_freq_anemometre_new_signal : in  std_logic                    := '0';             -- anemometer_in_freq_anemometre.new_signal
		clk_clk                                  : in  std_logic                    := '0';             --                           clk.clk
		keys_in_export                           : in  std_logic_vector(1 downto 0) := (others => '0'); --                       keys_in.export
		leds_out_export                          : out std_logic_vector(7 downto 0);                    --                      leds_out.export
		pwm_out_new_signal                       : out std_logic;                                       --                       pwm_out.new_signal
		reset_reset_n                            : in  std_logic                    := '0'              --                         reset.reset_n
	);
end entity SoC;

architecture rtl of SoC is
	component anemometre_avalon is
		port (
			address            : in  std_logic                     := 'X';             -- address
			writedata          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			readdata           : out std_logic_vector(31 downto 0);                    -- readdata
			write_n            : in  std_logic                     := 'X';             -- write_n
			chipselect         : in  std_logic                     := 'X';             -- chipselect
			reset_n            : in  std_logic                     := 'X';             -- reset_n
			clk_50M            : in  std_logic                     := 'X';             -- clk
			in_freq_anemometre : in  std_logic                     := 'X';             -- new_signal
			data_anemometre    : out std_logic_vector(7 downto 0);                     -- new_signal
			data_valid         : out std_logic                                         -- new_signal
		);
	end component anemometre_avalon;

	component SoC_KEYs is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(1 downto 0)  := (others => 'X')  -- export
		);
	end component SoC_KEYs;

	component SoC_LEDs is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(7 downto 0)                      -- export
		);
	end component SoC_LEDs;

	component SoC_NIOS_MCU is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(17 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(17 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component SoC_NIOS_MCU;

	component pwm_avalon is
		generic (
			freq_bus : integer := 16;
			duty_bus : integer := 16
		);
		port (
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			write_n    : in  std_logic                     := 'X';             -- write_n
			chipselect : in  std_logic                     := 'X';             -- chipselect
			clock      : in  std_logic                     := 'X';             -- clk
			pwm_out    : out std_logic                                         -- new_signal
		);
	end component pwm_avalon;

	component SoC_SRAM is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(13 downto 0) := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X';             -- reset_req
			freeze     : in  std_logic                     := 'X'              -- freeze
		);
	end component SoC_SRAM;

	component SoC_jtag is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component SoC_jtag;

	component SoC_mm_interconnect_0 is
		port (
			clk_0_clk_clk                              : in  std_logic                     := 'X';             -- clk
			NIOS_MCU_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			PWM_reset_reset_bridge_in_reset_reset      : in  std_logic                     := 'X';             -- reset
			NIOS_MCU_data_master_address               : in  std_logic_vector(17 downto 0) := (others => 'X'); -- address
			NIOS_MCU_data_master_waitrequest           : out std_logic;                                        -- waitrequest
			NIOS_MCU_data_master_byteenable            : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			NIOS_MCU_data_master_read                  : in  std_logic                     := 'X';             -- read
			NIOS_MCU_data_master_readdata              : out std_logic_vector(31 downto 0);                    -- readdata
			NIOS_MCU_data_master_write                 : in  std_logic                     := 'X';             -- write
			NIOS_MCU_data_master_writedata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			NIOS_MCU_data_master_debugaccess           : in  std_logic                     := 'X';             -- debugaccess
			NIOS_MCU_instruction_master_address        : in  std_logic_vector(17 downto 0) := (others => 'X'); -- address
			NIOS_MCU_instruction_master_waitrequest    : out std_logic;                                        -- waitrequest
			NIOS_MCU_instruction_master_read           : in  std_logic                     := 'X';             -- read
			NIOS_MCU_instruction_master_readdata       : out std_logic_vector(31 downto 0);                    -- readdata
			Anemometer_avalon_slave_0_address          : out std_logic_vector(0 downto 0);                     -- address
			Anemometer_avalon_slave_0_write            : out std_logic;                                        -- write
			Anemometer_avalon_slave_0_readdata         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			Anemometer_avalon_slave_0_writedata        : out std_logic_vector(31 downto 0);                    -- writedata
			Anemometer_avalon_slave_0_chipselect       : out std_logic;                                        -- chipselect
			jtag_avalon_jtag_slave_address             : out std_logic_vector(0 downto 0);                     -- address
			jtag_avalon_jtag_slave_write               : out std_logic;                                        -- write
			jtag_avalon_jtag_slave_read                : out std_logic;                                        -- read
			jtag_avalon_jtag_slave_readdata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			jtag_avalon_jtag_slave_writedata           : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_avalon_jtag_slave_waitrequest         : in  std_logic                     := 'X';             -- waitrequest
			jtag_avalon_jtag_slave_chipselect          : out std_logic;                                        -- chipselect
			KEYs_s1_address                            : out std_logic_vector(1 downto 0);                     -- address
			KEYs_s1_readdata                           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			LEDs_s1_address                            : out std_logic_vector(1 downto 0);                     -- address
			LEDs_s1_write                              : out std_logic;                                        -- write
			LEDs_s1_readdata                           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			LEDs_s1_writedata                          : out std_logic_vector(31 downto 0);                    -- writedata
			LEDs_s1_chipselect                         : out std_logic;                                        -- chipselect
			NIOS_MCU_debug_mem_slave_address           : out std_logic_vector(8 downto 0);                     -- address
			NIOS_MCU_debug_mem_slave_write             : out std_logic;                                        -- write
			NIOS_MCU_debug_mem_slave_read              : out std_logic;                                        -- read
			NIOS_MCU_debug_mem_slave_readdata          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			NIOS_MCU_debug_mem_slave_writedata         : out std_logic_vector(31 downto 0);                    -- writedata
			NIOS_MCU_debug_mem_slave_byteenable        : out std_logic_vector(3 downto 0);                     -- byteenable
			NIOS_MCU_debug_mem_slave_waitrequest       : in  std_logic                     := 'X';             -- waitrequest
			NIOS_MCU_debug_mem_slave_debugaccess       : out std_logic;                                        -- debugaccess
			PWM_avalon_slave_0_address                 : out std_logic_vector(1 downto 0);                     -- address
			PWM_avalon_slave_0_write                   : out std_logic;                                        -- write
			PWM_avalon_slave_0_readdata                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			PWM_avalon_slave_0_writedata               : out std_logic_vector(31 downto 0);                    -- writedata
			PWM_avalon_slave_0_chipselect              : out std_logic;                                        -- chipselect
			SRAM_s1_address                            : out std_logic_vector(13 downto 0);                    -- address
			SRAM_s1_write                              : out std_logic;                                        -- write
			SRAM_s1_readdata                           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			SRAM_s1_writedata                          : out std_logic_vector(31 downto 0);                    -- writedata
			SRAM_s1_byteenable                         : out std_logic_vector(3 downto 0);                     -- byteenable
			SRAM_s1_chipselect                         : out std_logic;                                        -- chipselect
			SRAM_s1_clken                              : out std_logic                                         -- clken
		);
	end component SoC_mm_interconnect_0;

	component SoC_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component SoC_irq_mapper;

	component soc_rst_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_in1      : in  std_logic := 'X';
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req      : out std_logic;
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component soc_rst_controller;

	component soc_rst_controller_001 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			reset_in1      : in  std_logic := 'X'; -- reset_in1.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_req      : out std_logic;        --          .reset_req
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component soc_rst_controller_001;

	signal nios_mcu_data_master_readdata                               : std_logic_vector(31 downto 0); -- mm_interconnect_0:NIOS_MCU_data_master_readdata -> NIOS_MCU:d_readdata
	signal nios_mcu_data_master_waitrequest                            : std_logic;                     -- mm_interconnect_0:NIOS_MCU_data_master_waitrequest -> NIOS_MCU:d_waitrequest
	signal nios_mcu_data_master_debugaccess                            : std_logic;                     -- NIOS_MCU:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:NIOS_MCU_data_master_debugaccess
	signal nios_mcu_data_master_address                                : std_logic_vector(17 downto 0); -- NIOS_MCU:d_address -> mm_interconnect_0:NIOS_MCU_data_master_address
	signal nios_mcu_data_master_byteenable                             : std_logic_vector(3 downto 0);  -- NIOS_MCU:d_byteenable -> mm_interconnect_0:NIOS_MCU_data_master_byteenable
	signal nios_mcu_data_master_read                                   : std_logic;                     -- NIOS_MCU:d_read -> mm_interconnect_0:NIOS_MCU_data_master_read
	signal nios_mcu_data_master_write                                  : std_logic;                     -- NIOS_MCU:d_write -> mm_interconnect_0:NIOS_MCU_data_master_write
	signal nios_mcu_data_master_writedata                              : std_logic_vector(31 downto 0); -- NIOS_MCU:d_writedata -> mm_interconnect_0:NIOS_MCU_data_master_writedata
	signal nios_mcu_instruction_master_readdata                        : std_logic_vector(31 downto 0); -- mm_interconnect_0:NIOS_MCU_instruction_master_readdata -> NIOS_MCU:i_readdata
	signal nios_mcu_instruction_master_waitrequest                     : std_logic;                     -- mm_interconnect_0:NIOS_MCU_instruction_master_waitrequest -> NIOS_MCU:i_waitrequest
	signal nios_mcu_instruction_master_address                         : std_logic_vector(17 downto 0); -- NIOS_MCU:i_address -> mm_interconnect_0:NIOS_MCU_instruction_master_address
	signal nios_mcu_instruction_master_read                            : std_logic;                     -- NIOS_MCU:i_read -> mm_interconnect_0:NIOS_MCU_instruction_master_read
	signal mm_interconnect_0_jtag_avalon_jtag_slave_chipselect         : std_logic;                     -- mm_interconnect_0:jtag_avalon_jtag_slave_chipselect -> jtag:av_chipselect
	signal mm_interconnect_0_jtag_avalon_jtag_slave_readdata           : std_logic_vector(31 downto 0); -- jtag:av_readdata -> mm_interconnect_0:jtag_avalon_jtag_slave_readdata
	signal mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest        : std_logic;                     -- jtag:av_waitrequest -> mm_interconnect_0:jtag_avalon_jtag_slave_waitrequest
	signal mm_interconnect_0_jtag_avalon_jtag_slave_address            : std_logic_vector(0 downto 0);  -- mm_interconnect_0:jtag_avalon_jtag_slave_address -> jtag:av_address
	signal mm_interconnect_0_jtag_avalon_jtag_slave_read               : std_logic;                     -- mm_interconnect_0:jtag_avalon_jtag_slave_read -> mm_interconnect_0_jtag_avalon_jtag_slave_read:in
	signal mm_interconnect_0_jtag_avalon_jtag_slave_write              : std_logic;                     -- mm_interconnect_0:jtag_avalon_jtag_slave_write -> mm_interconnect_0_jtag_avalon_jtag_slave_write:in
	signal mm_interconnect_0_jtag_avalon_jtag_slave_writedata          : std_logic_vector(31 downto 0); -- mm_interconnect_0:jtag_avalon_jtag_slave_writedata -> jtag:av_writedata
	signal mm_interconnect_0_pwm_avalon_slave_0_chipselect             : std_logic;                     -- mm_interconnect_0:PWM_avalon_slave_0_chipselect -> PWM:chipselect
	signal mm_interconnect_0_pwm_avalon_slave_0_readdata               : std_logic_vector(31 downto 0); -- PWM:readdata -> mm_interconnect_0:PWM_avalon_slave_0_readdata
	signal mm_interconnect_0_pwm_avalon_slave_0_address                : std_logic_vector(1 downto 0);  -- mm_interconnect_0:PWM_avalon_slave_0_address -> PWM:address
	signal mm_interconnect_0_pwm_avalon_slave_0_write                  : std_logic;                     -- mm_interconnect_0:PWM_avalon_slave_0_write -> mm_interconnect_0_pwm_avalon_slave_0_write:in
	signal mm_interconnect_0_pwm_avalon_slave_0_writedata              : std_logic_vector(31 downto 0); -- mm_interconnect_0:PWM_avalon_slave_0_writedata -> PWM:writedata
	signal mm_interconnect_0_anemometer_avalon_slave_0_chipselect      : std_logic;                     -- mm_interconnect_0:Anemometer_avalon_slave_0_chipselect -> Anemometer:chipselect
	signal mm_interconnect_0_anemometer_avalon_slave_0_readdata        : std_logic_vector(31 downto 0); -- Anemometer:readdata -> mm_interconnect_0:Anemometer_avalon_slave_0_readdata
	signal mm_interconnect_0_anemometer_avalon_slave_0_address         : std_logic_vector(0 downto 0);  -- mm_interconnect_0:Anemometer_avalon_slave_0_address -> Anemometer:address
	signal mm_interconnect_0_anemometer_avalon_slave_0_write           : std_logic;                     -- mm_interconnect_0:Anemometer_avalon_slave_0_write -> mm_interconnect_0_anemometer_avalon_slave_0_write:in
	signal mm_interconnect_0_anemometer_avalon_slave_0_writedata       : std_logic_vector(31 downto 0); -- mm_interconnect_0:Anemometer_avalon_slave_0_writedata -> Anemometer:writedata
	signal mm_interconnect_0_nios_mcu_debug_mem_slave_readdata         : std_logic_vector(31 downto 0); -- NIOS_MCU:debug_mem_slave_readdata -> mm_interconnect_0:NIOS_MCU_debug_mem_slave_readdata
	signal mm_interconnect_0_nios_mcu_debug_mem_slave_waitrequest      : std_logic;                     -- NIOS_MCU:debug_mem_slave_waitrequest -> mm_interconnect_0:NIOS_MCU_debug_mem_slave_waitrequest
	signal mm_interconnect_0_nios_mcu_debug_mem_slave_debugaccess      : std_logic;                     -- mm_interconnect_0:NIOS_MCU_debug_mem_slave_debugaccess -> NIOS_MCU:debug_mem_slave_debugaccess
	signal mm_interconnect_0_nios_mcu_debug_mem_slave_address          : std_logic_vector(8 downto 0);  -- mm_interconnect_0:NIOS_MCU_debug_mem_slave_address -> NIOS_MCU:debug_mem_slave_address
	signal mm_interconnect_0_nios_mcu_debug_mem_slave_read             : std_logic;                     -- mm_interconnect_0:NIOS_MCU_debug_mem_slave_read -> NIOS_MCU:debug_mem_slave_read
	signal mm_interconnect_0_nios_mcu_debug_mem_slave_byteenable       : std_logic_vector(3 downto 0);  -- mm_interconnect_0:NIOS_MCU_debug_mem_slave_byteenable -> NIOS_MCU:debug_mem_slave_byteenable
	signal mm_interconnect_0_nios_mcu_debug_mem_slave_write            : std_logic;                     -- mm_interconnect_0:NIOS_MCU_debug_mem_slave_write -> NIOS_MCU:debug_mem_slave_write
	signal mm_interconnect_0_nios_mcu_debug_mem_slave_writedata        : std_logic_vector(31 downto 0); -- mm_interconnect_0:NIOS_MCU_debug_mem_slave_writedata -> NIOS_MCU:debug_mem_slave_writedata
	signal mm_interconnect_0_sram_s1_chipselect                        : std_logic;                     -- mm_interconnect_0:SRAM_s1_chipselect -> SRAM:chipselect
	signal mm_interconnect_0_sram_s1_readdata                          : std_logic_vector(31 downto 0); -- SRAM:readdata -> mm_interconnect_0:SRAM_s1_readdata
	signal mm_interconnect_0_sram_s1_address                           : std_logic_vector(13 downto 0); -- mm_interconnect_0:SRAM_s1_address -> SRAM:address
	signal mm_interconnect_0_sram_s1_byteenable                        : std_logic_vector(3 downto 0);  -- mm_interconnect_0:SRAM_s1_byteenable -> SRAM:byteenable
	signal mm_interconnect_0_sram_s1_write                             : std_logic;                     -- mm_interconnect_0:SRAM_s1_write -> SRAM:write
	signal mm_interconnect_0_sram_s1_writedata                         : std_logic_vector(31 downto 0); -- mm_interconnect_0:SRAM_s1_writedata -> SRAM:writedata
	signal mm_interconnect_0_sram_s1_clken                             : std_logic;                     -- mm_interconnect_0:SRAM_s1_clken -> SRAM:clken
	signal mm_interconnect_0_leds_s1_chipselect                        : std_logic;                     -- mm_interconnect_0:LEDs_s1_chipselect -> LEDs:chipselect
	signal mm_interconnect_0_leds_s1_readdata                          : std_logic_vector(31 downto 0); -- LEDs:readdata -> mm_interconnect_0:LEDs_s1_readdata
	signal mm_interconnect_0_leds_s1_address                           : std_logic_vector(1 downto 0);  -- mm_interconnect_0:LEDs_s1_address -> LEDs:address
	signal mm_interconnect_0_leds_s1_write                             : std_logic;                     -- mm_interconnect_0:LEDs_s1_write -> mm_interconnect_0_leds_s1_write:in
	signal mm_interconnect_0_leds_s1_writedata                         : std_logic_vector(31 downto 0); -- mm_interconnect_0:LEDs_s1_writedata -> LEDs:writedata
	signal mm_interconnect_0_keys_s1_readdata                          : std_logic_vector(31 downto 0); -- KEYs:readdata -> mm_interconnect_0:KEYs_s1_readdata
	signal mm_interconnect_0_keys_s1_address                           : std_logic_vector(1 downto 0);  -- mm_interconnect_0:KEYs_s1_address -> KEYs:address
	signal irq_mapper_receiver0_irq                                    : std_logic;                     -- jtag:av_irq -> irq_mapper:receiver0_irq
	signal nios_mcu_irq_irq                                            : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> NIOS_MCU:irq
	signal rst_controller_reset_out_reset                              : std_logic;                     -- rst_controller:reset_out -> [mm_interconnect_0:PWM_reset_reset_bridge_in_reset_reset, rst_controller_reset_out_reset:in]
	signal rst_controller_001_reset_out_reset                          : std_logic;                     -- rst_controller_001:reset_out -> [SRAM:reset, irq_mapper:reset, mm_interconnect_0:NIOS_MCU_reset_reset_bridge_in_reset_reset, rst_controller_001_reset_out_reset:in, rst_translator:in_reset]
	signal rst_controller_001_reset_out_reset_req                      : std_logic;                     -- rst_controller_001:reset_req -> [NIOS_MCU:reset_req, SRAM:reset_req, rst_translator:reset_req_in]
	signal nios_mcu_debug_reset_request_reset                          : std_logic;                     -- NIOS_MCU:debug_reset_request -> rst_controller_001:reset_in1
	signal reset_reset_n_ports_inv                                     : std_logic;                     -- reset_reset_n:inv -> [rst_controller:reset_in0, rst_controller_001:reset_in0]
	signal mm_interconnect_0_jtag_avalon_jtag_slave_read_ports_inv     : std_logic;                     -- mm_interconnect_0_jtag_avalon_jtag_slave_read:inv -> jtag:av_read_n
	signal mm_interconnect_0_jtag_avalon_jtag_slave_write_ports_inv    : std_logic;                     -- mm_interconnect_0_jtag_avalon_jtag_slave_write:inv -> jtag:av_write_n
	signal mm_interconnect_0_pwm_avalon_slave_0_write_ports_inv        : std_logic;                     -- mm_interconnect_0_pwm_avalon_slave_0_write:inv -> PWM:write_n
	signal mm_interconnect_0_anemometer_avalon_slave_0_write_ports_inv : std_logic;                     -- mm_interconnect_0_anemometer_avalon_slave_0_write:inv -> Anemometer:write_n
	signal mm_interconnect_0_leds_s1_write_ports_inv                   : std_logic;                     -- mm_interconnect_0_leds_s1_write:inv -> LEDs:write_n
	signal rst_controller_reset_out_reset_ports_inv                    : std_logic;                     -- rst_controller_reset_out_reset:inv -> [Anemometer:reset_n, KEYs:reset_n, LEDs:reset_n, PWM:reset_n]
	signal rst_controller_001_reset_out_reset_ports_inv                : std_logic;                     -- rst_controller_001_reset_out_reset:inv -> [NIOS_MCU:reset_n, jtag:rst_n]

begin

	anemometer : component anemometre_avalon
		port map (
			address            => mm_interconnect_0_anemometer_avalon_slave_0_address(0),      --     avalon_slave_0.address
			writedata          => mm_interconnect_0_anemometer_avalon_slave_0_writedata,       --                   .writedata
			readdata           => mm_interconnect_0_anemometer_avalon_slave_0_readdata,        --                   .readdata
			write_n            => mm_interconnect_0_anemometer_avalon_slave_0_write_ports_inv, --                   .write_n
			chipselect         => mm_interconnect_0_anemometer_avalon_slave_0_chipselect,      --                   .chipselect
			reset_n            => rst_controller_reset_out_reset_ports_inv,                    --              reset.reset_n
			clk_50M            => clk_clk,                                                     --              clock.clk
			in_freq_anemometre => anemometer_in_freq_anemometre_new_signal,                    -- in_freq_anemometre.new_signal
			data_anemometre    => anemometer_data_anemometre_new_signal,                       --    data_anemometre.new_signal
			data_valid         => anemometer_data_valid_new_signal                             --         data_valid.new_signal
		);

	keys : component SoC_KEYs
		port map (
			clk      => clk_clk,                                  --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv, --               reset.reset_n
			address  => mm_interconnect_0_keys_s1_address,        --                  s1.address
			readdata => mm_interconnect_0_keys_s1_readdata,       --                    .readdata
			in_port  => keys_in_export                            -- external_connection.export
		);

	leds : component SoC_LEDs
		port map (
			clk        => clk_clk,                                   --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,  --               reset.reset_n
			address    => mm_interconnect_0_leds_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_leds_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_leds_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_leds_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_leds_s1_readdata,        --                    .readdata
			out_port   => leds_out_export                            -- external_connection.export
		);

	nios_mcu : component SoC_NIOS_MCU
		port map (
			clk                                 => clk_clk,                                                --                       clk.clk
			reset_n                             => rst_controller_001_reset_out_reset_ports_inv,           --                     reset.reset_n
			reset_req                           => rst_controller_001_reset_out_reset_req,                 --                          .reset_req
			d_address                           => nios_mcu_data_master_address,                           --               data_master.address
			d_byteenable                        => nios_mcu_data_master_byteenable,                        --                          .byteenable
			d_read                              => nios_mcu_data_master_read,                              --                          .read
			d_readdata                          => nios_mcu_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => nios_mcu_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => nios_mcu_data_master_write,                             --                          .write
			d_writedata                         => nios_mcu_data_master_writedata,                         --                          .writedata
			debug_mem_slave_debugaccess_to_roms => nios_mcu_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => nios_mcu_instruction_master_address,                    --        instruction_master.address
			i_read                              => nios_mcu_instruction_master_read,                       --                          .read
			i_readdata                          => nios_mcu_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => nios_mcu_instruction_master_waitrequest,                --                          .waitrequest
			irq                                 => nios_mcu_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => nios_mcu_debug_reset_request_reset,                     --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_0_nios_mcu_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_0_nios_mcu_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_0_nios_mcu_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_0_nios_mcu_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_0_nios_mcu_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_0_nios_mcu_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_0_nios_mcu_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_0_nios_mcu_debug_mem_slave_writedata,   --                          .writedata
			dummy_ci_port                       => open                                                    -- custom_instruction_master.readra
		);

	pwm : component pwm_avalon
		generic map (
			freq_bus => 16,
			duty_bus => 16
		)
		port map (
			reset_n    => rst_controller_reset_out_reset_ports_inv,             --          reset.reset_n
			address    => mm_interconnect_0_pwm_avalon_slave_0_address,         -- avalon_slave_0.address
			writedata  => mm_interconnect_0_pwm_avalon_slave_0_writedata,       --               .writedata
			readdata   => mm_interconnect_0_pwm_avalon_slave_0_readdata,        --               .readdata
			write_n    => mm_interconnect_0_pwm_avalon_slave_0_write_ports_inv, --               .write_n
			chipselect => mm_interconnect_0_pwm_avalon_slave_0_chipselect,      --               .chipselect
			clock      => clk_clk,                                              --          clock.clk
			pwm_out    => pwm_out_new_signal                                    --        pwm_out.new_signal
		);

	sram : component SoC_SRAM
		port map (
			clk        => clk_clk,                                --   clk1.clk
			address    => mm_interconnect_0_sram_s1_address,      --     s1.address
			clken      => mm_interconnect_0_sram_s1_clken,        --       .clken
			chipselect => mm_interconnect_0_sram_s1_chipselect,   --       .chipselect
			write      => mm_interconnect_0_sram_s1_write,        --       .write
			readdata   => mm_interconnect_0_sram_s1_readdata,     --       .readdata
			writedata  => mm_interconnect_0_sram_s1_writedata,    --       .writedata
			byteenable => mm_interconnect_0_sram_s1_byteenable,   --       .byteenable
			reset      => rst_controller_001_reset_out_reset,     -- reset1.reset
			reset_req  => rst_controller_001_reset_out_reset_req, --       .reset_req
			freeze     => '0'                                     -- (terminated)
		);

	jtag : component SoC_jtag
		port map (
			clk            => clk_clk,                                                  --               clk.clk
			rst_n          => rst_controller_001_reset_out_reset_ports_inv,             --             reset.reset_n
			av_chipselect  => mm_interconnect_0_jtag_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_0_jtag_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_0_jtag_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_0_jtag_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_0_jtag_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_0_jtag_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver0_irq                                  --               irq.irq
		);

	mm_interconnect_0 : component SoC_mm_interconnect_0
		port map (
			clk_0_clk_clk                              => clk_clk,                                                --                            clk_0_clk.clk
			NIOS_MCU_reset_reset_bridge_in_reset_reset => rst_controller_001_reset_out_reset,                     -- NIOS_MCU_reset_reset_bridge_in_reset.reset
			PWM_reset_reset_bridge_in_reset_reset      => rst_controller_reset_out_reset,                         --      PWM_reset_reset_bridge_in_reset.reset
			NIOS_MCU_data_master_address               => nios_mcu_data_master_address,                           --                 NIOS_MCU_data_master.address
			NIOS_MCU_data_master_waitrequest           => nios_mcu_data_master_waitrequest,                       --                                     .waitrequest
			NIOS_MCU_data_master_byteenable            => nios_mcu_data_master_byteenable,                        --                                     .byteenable
			NIOS_MCU_data_master_read                  => nios_mcu_data_master_read,                              --                                     .read
			NIOS_MCU_data_master_readdata              => nios_mcu_data_master_readdata,                          --                                     .readdata
			NIOS_MCU_data_master_write                 => nios_mcu_data_master_write,                             --                                     .write
			NIOS_MCU_data_master_writedata             => nios_mcu_data_master_writedata,                         --                                     .writedata
			NIOS_MCU_data_master_debugaccess           => nios_mcu_data_master_debugaccess,                       --                                     .debugaccess
			NIOS_MCU_instruction_master_address        => nios_mcu_instruction_master_address,                    --          NIOS_MCU_instruction_master.address
			NIOS_MCU_instruction_master_waitrequest    => nios_mcu_instruction_master_waitrequest,                --                                     .waitrequest
			NIOS_MCU_instruction_master_read           => nios_mcu_instruction_master_read,                       --                                     .read
			NIOS_MCU_instruction_master_readdata       => nios_mcu_instruction_master_readdata,                   --                                     .readdata
			Anemometer_avalon_slave_0_address          => mm_interconnect_0_anemometer_avalon_slave_0_address,    --            Anemometer_avalon_slave_0.address
			Anemometer_avalon_slave_0_write            => mm_interconnect_0_anemometer_avalon_slave_0_write,      --                                     .write
			Anemometer_avalon_slave_0_readdata         => mm_interconnect_0_anemometer_avalon_slave_0_readdata,   --                                     .readdata
			Anemometer_avalon_slave_0_writedata        => mm_interconnect_0_anemometer_avalon_slave_0_writedata,  --                                     .writedata
			Anemometer_avalon_slave_0_chipselect       => mm_interconnect_0_anemometer_avalon_slave_0_chipselect, --                                     .chipselect
			jtag_avalon_jtag_slave_address             => mm_interconnect_0_jtag_avalon_jtag_slave_address,       --               jtag_avalon_jtag_slave.address
			jtag_avalon_jtag_slave_write               => mm_interconnect_0_jtag_avalon_jtag_slave_write,         --                                     .write
			jtag_avalon_jtag_slave_read                => mm_interconnect_0_jtag_avalon_jtag_slave_read,          --                                     .read
			jtag_avalon_jtag_slave_readdata            => mm_interconnect_0_jtag_avalon_jtag_slave_readdata,      --                                     .readdata
			jtag_avalon_jtag_slave_writedata           => mm_interconnect_0_jtag_avalon_jtag_slave_writedata,     --                                     .writedata
			jtag_avalon_jtag_slave_waitrequest         => mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest,   --                                     .waitrequest
			jtag_avalon_jtag_slave_chipselect          => mm_interconnect_0_jtag_avalon_jtag_slave_chipselect,    --                                     .chipselect
			KEYs_s1_address                            => mm_interconnect_0_keys_s1_address,                      --                              KEYs_s1.address
			KEYs_s1_readdata                           => mm_interconnect_0_keys_s1_readdata,                     --                                     .readdata
			LEDs_s1_address                            => mm_interconnect_0_leds_s1_address,                      --                              LEDs_s1.address
			LEDs_s1_write                              => mm_interconnect_0_leds_s1_write,                        --                                     .write
			LEDs_s1_readdata                           => mm_interconnect_0_leds_s1_readdata,                     --                                     .readdata
			LEDs_s1_writedata                          => mm_interconnect_0_leds_s1_writedata,                    --                                     .writedata
			LEDs_s1_chipselect                         => mm_interconnect_0_leds_s1_chipselect,                   --                                     .chipselect
			NIOS_MCU_debug_mem_slave_address           => mm_interconnect_0_nios_mcu_debug_mem_slave_address,     --             NIOS_MCU_debug_mem_slave.address
			NIOS_MCU_debug_mem_slave_write             => mm_interconnect_0_nios_mcu_debug_mem_slave_write,       --                                     .write
			NIOS_MCU_debug_mem_slave_read              => mm_interconnect_0_nios_mcu_debug_mem_slave_read,        --                                     .read
			NIOS_MCU_debug_mem_slave_readdata          => mm_interconnect_0_nios_mcu_debug_mem_slave_readdata,    --                                     .readdata
			NIOS_MCU_debug_mem_slave_writedata         => mm_interconnect_0_nios_mcu_debug_mem_slave_writedata,   --                                     .writedata
			NIOS_MCU_debug_mem_slave_byteenable        => mm_interconnect_0_nios_mcu_debug_mem_slave_byteenable,  --                                     .byteenable
			NIOS_MCU_debug_mem_slave_waitrequest       => mm_interconnect_0_nios_mcu_debug_mem_slave_waitrequest, --                                     .waitrequest
			NIOS_MCU_debug_mem_slave_debugaccess       => mm_interconnect_0_nios_mcu_debug_mem_slave_debugaccess, --                                     .debugaccess
			PWM_avalon_slave_0_address                 => mm_interconnect_0_pwm_avalon_slave_0_address,           --                   PWM_avalon_slave_0.address
			PWM_avalon_slave_0_write                   => mm_interconnect_0_pwm_avalon_slave_0_write,             --                                     .write
			PWM_avalon_slave_0_readdata                => mm_interconnect_0_pwm_avalon_slave_0_readdata,          --                                     .readdata
			PWM_avalon_slave_0_writedata               => mm_interconnect_0_pwm_avalon_slave_0_writedata,         --                                     .writedata
			PWM_avalon_slave_0_chipselect              => mm_interconnect_0_pwm_avalon_slave_0_chipselect,        --                                     .chipselect
			SRAM_s1_address                            => mm_interconnect_0_sram_s1_address,                      --                              SRAM_s1.address
			SRAM_s1_write                              => mm_interconnect_0_sram_s1_write,                        --                                     .write
			SRAM_s1_readdata                           => mm_interconnect_0_sram_s1_readdata,                     --                                     .readdata
			SRAM_s1_writedata                          => mm_interconnect_0_sram_s1_writedata,                    --                                     .writedata
			SRAM_s1_byteenable                         => mm_interconnect_0_sram_s1_byteenable,                   --                                     .byteenable
			SRAM_s1_chipselect                         => mm_interconnect_0_sram_s1_chipselect,                   --                                     .chipselect
			SRAM_s1_clken                              => mm_interconnect_0_sram_s1_clken                         --                                     .clken
		);

	irq_mapper : component SoC_irq_mapper
		port map (
			clk           => clk_clk,                            --       clk.clk
			reset         => rst_controller_001_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,           -- receiver0.irq
			sender_irq    => nios_mcu_irq_irq                    --    sender.irq
		);

	rst_controller : component soc_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,        -- reset_in0.reset
			clk            => clk_clk,                        --       clk.clk
			reset_out      => rst_controller_reset_out_reset, -- reset_out.reset
			reset_req      => open,                           -- (terminated)
			reset_req_in0  => '0',                            -- (terminated)
			reset_in1      => '0',                            -- (terminated)
			reset_req_in1  => '0',                            -- (terminated)
			reset_in2      => '0',                            -- (terminated)
			reset_req_in2  => '0',                            -- (terminated)
			reset_in3      => '0',                            -- (terminated)
			reset_req_in3  => '0',                            -- (terminated)
			reset_in4      => '0',                            -- (terminated)
			reset_req_in4  => '0',                            -- (terminated)
			reset_in5      => '0',                            -- (terminated)
			reset_req_in5  => '0',                            -- (terminated)
			reset_in6      => '0',                            -- (terminated)
			reset_req_in6  => '0',                            -- (terminated)
			reset_in7      => '0',                            -- (terminated)
			reset_req_in7  => '0',                            -- (terminated)
			reset_in8      => '0',                            -- (terminated)
			reset_req_in8  => '0',                            -- (terminated)
			reset_in9      => '0',                            -- (terminated)
			reset_req_in9  => '0',                            -- (terminated)
			reset_in10     => '0',                            -- (terminated)
			reset_req_in10 => '0',                            -- (terminated)
			reset_in11     => '0',                            -- (terminated)
			reset_req_in11 => '0',                            -- (terminated)
			reset_in12     => '0',                            -- (terminated)
			reset_req_in12 => '0',                            -- (terminated)
			reset_in13     => '0',                            -- (terminated)
			reset_req_in13 => '0',                            -- (terminated)
			reset_in14     => '0',                            -- (terminated)
			reset_req_in14 => '0',                            -- (terminated)
			reset_in15     => '0',                            -- (terminated)
			reset_req_in15 => '0'                             -- (terminated)
		);

	rst_controller_001 : component soc_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,                -- reset_in0.reset
			reset_in1      => nios_mcu_debug_reset_request_reset,     -- reset_in1.reset
			clk            => clk_clk,                                --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_001_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                    -- (terminated)
			reset_req_in1  => '0',                                    -- (terminated)
			reset_in2      => '0',                                    -- (terminated)
			reset_req_in2  => '0',                                    -- (terminated)
			reset_in3      => '0',                                    -- (terminated)
			reset_req_in3  => '0',                                    -- (terminated)
			reset_in4      => '0',                                    -- (terminated)
			reset_req_in4  => '0',                                    -- (terminated)
			reset_in5      => '0',                                    -- (terminated)
			reset_req_in5  => '0',                                    -- (terminated)
			reset_in6      => '0',                                    -- (terminated)
			reset_req_in6  => '0',                                    -- (terminated)
			reset_in7      => '0',                                    -- (terminated)
			reset_req_in7  => '0',                                    -- (terminated)
			reset_in8      => '0',                                    -- (terminated)
			reset_req_in8  => '0',                                    -- (terminated)
			reset_in9      => '0',                                    -- (terminated)
			reset_req_in9  => '0',                                    -- (terminated)
			reset_in10     => '0',                                    -- (terminated)
			reset_req_in10 => '0',                                    -- (terminated)
			reset_in11     => '0',                                    -- (terminated)
			reset_req_in11 => '0',                                    -- (terminated)
			reset_in12     => '0',                                    -- (terminated)
			reset_req_in12 => '0',                                    -- (terminated)
			reset_in13     => '0',                                    -- (terminated)
			reset_req_in13 => '0',                                    -- (terminated)
			reset_in14     => '0',                                    -- (terminated)
			reset_req_in14 => '0',                                    -- (terminated)
			reset_in15     => '0',                                    -- (terminated)
			reset_req_in15 => '0'                                     -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	mm_interconnect_0_jtag_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_jtag_avalon_jtag_slave_read;

	mm_interconnect_0_jtag_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_jtag_avalon_jtag_slave_write;

	mm_interconnect_0_pwm_avalon_slave_0_write_ports_inv <= not mm_interconnect_0_pwm_avalon_slave_0_write;

	mm_interconnect_0_anemometer_avalon_slave_0_write_ports_inv <= not mm_interconnect_0_anemometer_avalon_slave_0_write;

	mm_interconnect_0_leds_s1_write_ports_inv <= not mm_interconnect_0_leds_s1_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

	rst_controller_001_reset_out_reset_ports_inv <= not rst_controller_001_reset_out_reset;

end architecture rtl; -- of SoC
